package tb_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
//`include "axi_if.sv"
`include "axi_trans.sv"
`include "axi_seq.sv"
`include "axi_sequencer.sv"
`include "axi_driver.sv"
`include "axi_monitor.sv"
`include "axi_coverage.sv"
`include "axi_agent.sv"
`include "axi_scoreboard.sv"
`include "axi_env.sv"
`include "test.sv"
endpackage
