class axi_agent extends uvm_agent;
  `uvm_component_utils(axi_agent)
  axi_driver driver;
  axi_monitor monitor;
  axi_sequencer sequencer;

  function new(string name = "axi_agent",uvm_component parent = null);
   super.new(name,parent);
   
  endfunction

  virtual function void build_phase(uvm_phase phase);
   super.build_phase(phase);
   driver = axi_driver::type_id::create("driver",this);  
   monitor = axi_monitor::type_id::create("monitor",this);  
   sequencer = axi_sequencer::type_id::create("sequencer",this);  
  endfunction

  virtual function void connect_phase(uvm_phase phase);
   if(get_is_active() == UVM_ACTIVE)
   begin
   driver.seq_item_port.connect(sequencer.seq_item_export);
   end
  endfunction
endclass
